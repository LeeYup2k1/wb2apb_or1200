
module 
endmodule
